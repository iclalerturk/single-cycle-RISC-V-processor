module instructionMemory(
    input [31:0] A,
    output reg [31:0] RD
    );
//wire [3:0] add = A[3:0];
reg [31:0] mem1[51:0];
initial begin
    mem1[0] = 32'b00000000011100110000001010110011; // add
    mem1[4] = 32'b01000000011100110000001010110011; // sub
    mem1[8] = 32'hFFC4A303; // lw 
    mem1[12] = 32'b11011110001110111101000011101111; //jal
    mem1[16] = 32'b11111111101100100010000110010011 ; // slti 
    mem1[20] = 32'hFE420AE3; // beq
    mem1[24] = 32'h0064A423; // sw
    mem1[28] = 32'b11111111111100110110001010010011; // ori 
    mem1[32] = 32'b00000000011100100000000110010011; // andi
    mem1[36] = 32'h0062E233; // or
    mem1[40] = 32'b00000000001000110000001010010011; // addi
    mem1[44] = 32'b00000000010100100010000110110011; // slt
    mem1[48] = 32'b00000000010100100111000110110011; // and


    
end
always @(*) begin
    RD = mem1[A]; 
end

endmodule